`define CLK_FREQ 50000000   // 50 MHz
`define BAUD_RATE 115200    // 11520 bytes/s ~ 11Kb/s
`define WIDTH 8             // one byte
